//Guia_0701.v
//Cauã Costa Alves

module Guia_0701 ( input a,
                   input b,
                   output op1,
                   output op2)